module DMA(
    // DMA Interface
    input wire  [15:0]  SRC,
    input wire  [15:0]  DST,
    input wire  [7:0]   LEN,
    input wire  [7:0]   INC,

    // INT Interface
    output wire INT_DONE,
    output wire INT_FAIL,

    output 
);


endmodule